BZh91AY&SYoq� u߀Px���g߰����P�9m��hРH��0��Ba4h�&�4 ɑ�i�j�)�       JdI��2��� P OS� �0# #	��14�H��0�M���1�4�� �DĒ{D�@��@H+	>���6���!���7�0@X4���چMX��6ݴD9P��m8LP�ƛ:ҭr�����jS��\�����RIӒ�'i���D�2����u�����./'���Az�L�.qh/d�$�E/H	C>ئ�D_��n*:-��/6�i�C�k��[�*E��g1�>Kl7���z�qY٦^ �|���C@ꈇ*�eKa@���:n혲q*3�(���H�W���A�<*�c�ʚj.����wV�&�8)Y�h��/$C�����������WR)�9�i;E�`��g(��,�f ND�jjL�����(R�S�*w�(�K�8cE�9br�A$��T�:��6��,W��#:��n�����^"��|g��>�1Ɛ���Q$�(�!����ƌ6���4w֓�ʫ�� $����Bf��AtQ�kR�0l�`뙭0���̧nG:f����W�I��<��G��?9H�L.Qen���ce���*���,V�W�!-j��bX���D��B_	�81��-��=`ʸD�!u���h�4+%�-���D3['�I P�-6�����D���[8"��R��WE�ՄБ�h�h	H�P�D��|e���-&V��&��6Q��P�1��+��!�N��)D�r��wb�1	F�1%{�*��)�YVAKsUh��<�<�1<O�2���=����t�a+Mx��	y��L[�+9d�4V��򳈣�H�s�O	\I&�Ā$�:�@�LL��N�9W"���<�%
a��b�uK���΢�{�,�@�v���WPC%������΃�٤$�$oLkg>b�$U3Q4�މ*�D�+D�H&;L�Y�U3�tޭ�W���_Y:����b��d8�-+HiȠcmu�7��1��a�Av�����S-�,3�h�]y���2T��ӕ�{�۫���"�(H7��׀